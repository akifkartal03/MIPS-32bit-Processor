module constant_producer(zero,one,two,three);
output [31:0] zero,one,two,three;


and a2(zero[0],0,1);
and a3(zero[1],0,1);
and a4(zero[2],0,1);
and a5(zero[3],0,1);
and a6(zero[4],0,1);
and a7(zero[5],0,1);
and a8(zero[6],0,1);
and a9(zero[7],0,1);
and a10(zero[8],0,1);
and a11(zero[9],0,1);
and a12(zero[10],0,1);
and a13(zero[11],0,1);
and a14(zero[12],0,1);
and a15(zero[13],0,1);
and a16(zero[14],0,1);
and a17(zero[15],0,1);
and a18(zero[16],0,1);
and a19(zero[17],0,1);
and a20(zero[18],0,1);
and a21(zero[19],0,1);
and a22(zero[20],0,1);
and a23(zero[21],0,1);
and a24(zero[22],0,1);
and a25(zero[23],0,1);
and a26(zero[24],0,1);
and a27(zero[25],0,1);
and a28(zero[26],0,1);
and a29(zero[27],0,1);
and a30(zero[28],0,1);
and a31(zero[29],0,1);
and a32(zero[30],0,1);
and a33(zero[31],0,1);


and a210(one[0],1,1);
and a311(one[1],0,1);
and a40(one[2],0,1);
and a50(one[3],0,1);
and a60(one[4],0,1);
and a70(one[5],0,1);
and a80(one[6],0,1);
and a90(one[7],0,1);
and a100(one[8],0,1);
and a110(one[9],0,1);
and a120(one[10],0,1);
and a130(one[11],0,1);
and a140(one[12],0,1);
and a150(one[13],0,1);
and a160(one[14],0,1);
and a170(one[15],0,1);
and a180(one[16],0,1);
and a190(one[17],0,1);
and a200(one[18],0,1);
and a2101(one[19],0,1);
and a220(one[20],0,1);
and a230(one[21],0,1);
and a240(one[22],0,1);
and a250(one[23],0,1);
and a260(one[24],0,1);
and a270(one[25],0,1);
and a280(one[26],0,1);
and a290(one[27],0,1);
and a300(one[28],0,1);
and a310(one[29],0,1);
and a320(one[30],0,1);
and a330(one[31],0,1);

and a289(two[0],0,1);
and a389(two[1],1,1);
and a41(two[2],0,1);
and a51(two[3],0,1);
and a61(two[4],0,1);
and a71(two[5],0,1);
and a81(two[6],0,1);
and a91(two[7],0,1);
and a101(two[8],0,1);
and a111(two[9],0,1);
and a121(two[10],0,1);
and a131(two[11],0,1);
and a141(two[12],0,1);
and a151(two[13],0,1);
and a161(two[14],0,1);
and a171(two[15],0,1);
and a181(two[16],0,1);
and a191(two[17],0,1);
and a201(two[18],0,1);
and a211(two[19],0,1);
and a221(two[20],0,1);
and a231(two[21],0,1);
and a241(two[22],0,1);
and a251(two[23],0,1);
and a261(two[24],0,1);
and a271(two[25],0,1);
and a281(two[26],0,1);
and a291(two[27],0,1);
and a301(two[28],0,1);
and a3111(two[29],0,1);
and a321(two[30],0,1);
and a331(two[31],0,1);

and a263(three[0],1,1);
and a369(three[1],1,1);
and a42(three[2],0,1);
and a52(three[3],0,1);
and a62(three[4],0,1);
and a72(three[5],0,1);
and a82(three[6],0,1);
and a92(three[7],0,1);
and a102(three[8],0,1);
and a112(three[9],0,1);
and a122(three[10],0,1);
and a132(three[11],0,1);
and a142(three[12],0,1);
and a152(three[13],0,1);
and a162(three[14],0,1);
and a172(three[15],0,1);
and a182(three[16],0,1);
and a192(three[17],0,1);
and a202(three[18],0,1);
and a212(three[19],0,1);
and a222(three[20],0,1);
and a232(three[21],0,1);
and a242(three[22],0,1);
and a252(three[23],0,1);
and a262(three[24],0,1);
and a272(three[25],0,1);
and a282(three[26],0,1);
and a292(three[27],0,1);
and a302(three[28],0,1);
and a312(three[29],0,1);
and a322(three[30],0,1);
and a332(three[31],0,1);

endmodule