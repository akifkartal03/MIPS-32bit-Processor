module alu_32bit_testbench();
	reg signed [31:0] a,b;
	reg [2:0] alu_ctr;
	wire c_out,z;
	wire signed [31:0] r;
	alu_32bit my_alu32(r,c_out,z,a,b,alu_ctr);
	initial begin
	//a=10, b=30
	a = 32'b00000000000000000000000000001010; b =32'b00000000000000000000000000011110; alu_ctr =3'b000; //and
	#20;
	//a=0, b=10
	a = 32'b00000000000000000000000000000000; b =32'b00000000000000000000000000010100; alu_ctr =3'b000; //and
	#20;
	//a=10, b=30
	a = 32'b00000000000000000000000000001010; b =32'b00000000000000000000000000011110; alu_ctr =3'b001; //or
	#20;
	//a=0, b=10
	a = 32'b00000000000000000000000000000000; b =32'b00000000000000000000000000010100; alu_ctr =3'b001; //or
	#20;
	//a=10, b=30
	a = 32'b00000000000000000000000000001010; b =32'b00000000000000000000000000011110; alu_ctr =3'b010; //add
	#20;
	//a=0, b=10
	a = 32'b00000000000000000000000000000000; b =32'b00000000000000000000000000010100; alu_ctr =3'b010; //add
	#20;
	//a=10, b=30
	a = 32'b00000000000000000000000000001010; b =32'b00000000000000000000000000011110; alu_ctr =3'b110; //sub
	#20;
	//a=0, b=10
	a = 32'b00000000000000000000000000000000; b =32'b00000000000000000000000000010100; alu_ctr =3'b110; //sub
	#20;
	//a=100, b=99
	a = 32'b00000000000000000000000001100100; b =32'b00000000000000000000000001100011; alu_ctr =3'b110; //sub
	#20;
	//a=10, b=30
	a = 32'b00000000000000000000000000001010; b =32'b00000000000000000000000000011110; alu_ctr =3'b111; //xor
	#20;
	//a=0, b=10
	a = 32'b00000000000000000000000000000000; b =32'b00000000000000000000000000010100; alu_ctr =3'b111; //xor
	#20;
	//a=10, b=10
	a = 32'b00000000000000000000000000010100; b =32'b00000000000000000000000000010100; alu_ctr =3'b111; //xor
	#20;
	end
	initial begin
	$monitor("time=%2d,a=%2d,b=%2d,alu_ctr=%3b,r=%2d,cout=%1b,z=%1b"
	          ,$time,a,b,alu_ctr,r,c_out,z);
	end
endmodule