module mux_32x1_testbench();
	reg [31:0] a;
	reg [31:0] b;
	wire [31:0] result;
	reg s0;
	mux_32x1 my_mux32(result,a,b,s0);
	initial begin
	a = 32'b00000_00000_00000_00000_00000_00000_00; b =32'b00000_00000_00000_00000_00000_01111_11; s0 = 1'b1;
	#20;
	a = 32'b00000_00000_00000_00000_00000_00000_00; b =32'b00000_00000_00000_00000_00000_01111_11; s0 = 1'b0;
	#20;
	a = 32'b00000_00000_00000_00100_00100_00100_10; b =32'b00000_00000_00000_00000_00000_01111_11; s0 = 1'b0;
	#20;
	end
	initial begin
	$monitor("time=%2d,a=%2d,b=%2d,s0=%1b,result=%2d",$time,a,b,s0,result);
	end
endmodule