module zero_extender(temp,number);
output [31:0] temp;
input [15:0] number;


and a2(temp[0],number[0],1);
and a3(temp[1],number[1],1);
and a4(temp[2],number[2],1);
and a5(temp[3],number[3],1);
and a6(temp[4],number[4],1);
and a7(temp[5],number[5],1);
and a8(temp[6],number[6],1);
and a9(temp[7],number[7],1);
and a10(temp[8],number[8],1);
and a11(temp[9],number[9],1);
and a12(temp[10],number[10],1);
and a13(temp[11],number[11],1);
and a14(temp[12],number[12],1);
and a15(temp[13],number[13],1);
and a16(temp[14],number[14],1);
and a17(temp[15],number[15],1);


and a18(temp[16],0,1);
and a19(temp[17],0,1);
and a20(temp[18],0,1);
and a21(temp[19],0,1);
and a22(temp[20],0,1);
and a23(temp[21],0,1);
and a24(temp[22],0,1);
and a25(temp[23],0,1);
and a26(temp[24],0,1);
and a27(temp[25],0,1);
and a28(temp[26],0,1);
and a29(temp[27],0,1);
and a30(temp[28],0,1);
and a31(temp[29],0,1);
and a32(temp[30],0,1);
and a33(temp[31],0,1);


endmodule