module mux_32x1(d,i0,i1,s0);
output [31:0] d;
input [31:0] i0,i1;
input s0;

mux_2x1 m1(d[0],i0[0],i1[0],s0);
mux_2x1 m2(d[1],i0[1],i1[1],s0);
mux_2x1 m3(d[2],i0[2],i1[2],s0);
mux_2x1 m4(d[3],i0[3],i1[3],s0);
mux_2x1 m5(d[4],i0[4],i1[4],s0);
mux_2x1 m6(d[5],i0[5],i1[5],s0);
mux_2x1 m7(d[6],i0[6],i1[6],s0);
mux_2x1 m8(d[7],i0[7],i1[7],s0);
mux_2x1 m9(d[8],i0[8],i1[8],s0);
mux_2x1 m10(d[9],i0[9],i1[9],s0);
mux_2x1 m11(d[10],i0[10],i1[10],s0);
mux_2x1 m12(d[11],i0[11],i1[11],s0);
mux_2x1 m13(d[12],i0[12],i1[12],s0);
mux_2x1 m14(d[13],i0[13],i1[13],s0);
mux_2x1 m15(d[14],i0[14],i1[14],s0);
mux_2x1 m16(d[15],i0[15],i1[15],s0);
mux_2x1 m17(d[16],i0[16],i1[16],s0);
mux_2x1 m18(d[17],i0[17],i1[17],s0);
mux_2x1 m19(d[18],i0[18],i1[18],s0);
mux_2x1 m20(d[19],i0[19],i1[19],s0);
mux_2x1 m21(d[20],i0[20],i1[20],s0);
mux_2x1 m22(d[21],i0[21],i1[21],s0);
mux_2x1 m23(d[22],i0[22],i1[22],s0);
mux_2x1 m24(d[23],i0[23],i1[23],s0);
mux_2x1 m25(d[24],i0[24],i1[24],s0);
mux_2x1 m26(d[25],i0[25],i1[25],s0);
mux_2x1 m27(d[26],i0[26],i1[26],s0);
mux_2x1 m28(d[27],i0[27],i1[27],s0);
mux_2x1 m29(d[28],i0[28],i1[28],s0);
mux_2x1 m30(d[29],i0[29],i1[29],s0);
mux_2x1 m31(d[30],i0[30],i1[30],s0);
mux_2x1 m32(d[31],i0[31],i1[31],s0);


endmodule